programa viko;
    var texto nombre;
realiza
    imprime("Cual es tu nombre?");
    lee(nombre);
    imprime("");
    imprime("Hola ",nombre,", esta es Sofi!");
fin
