programa jjj;
var numero x;
REALIZA
x = 10;
FIN

func numero uno(texto i)
realiza
  i = "hola";
fin
func numero dos(numero z, texto q)
var texto a;
realiza
a = "adios";
uno(a);
fin