programa viko;
    var numero i;
    var numero b;
    var numero a;
realiza
  para (i = 0; i mayor 8; i = i + 1;) realiza
    b = a + b;
  fin
fin