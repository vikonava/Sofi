programa viko;
var texto nombre
realiza
lee(nombre);
imprime("algo",nombre);
fin