programa viko;
    var numero c;
    var numero b;
    var numero a;
    var numero d;
realiza

a = 1;
b = 2 + 1;

fin