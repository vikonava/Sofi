programa viko;
    var booleano c;
    var numero b;
    var numero a;
realiza
  c = a mayor b;
fin