programa viko;
    var numero i;
    var numero j;
realiza
    para (j = 1; j menor 3; j = j + 1;) realiza
        para (i = 0; i menor 10; i = i + 1;) realiza
            imprime(i*j);
        fin
    fin
fin
