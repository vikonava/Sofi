programa viko;
    var numero nombre;
    var numero a;
realiza
    lee(nombre);
    imprime("algo",nombre); 
fin